** sch_path: /home/vlsi/Documents/sky130/inverter/xschem/pmos_char.sch
**.subckt pmos_char
Vgs g net1 0
XM1 net2 net1 g g sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vds g net2 0
Vds1 g GND 5
**** begin user architecture code
 .lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.dc Vds 0 1.8 1m Vgs 0 5 0.5
.save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
