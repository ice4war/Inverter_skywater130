magic
tech sky130A
timestamp 1706460133
<< nwell >>
rect -150 -100 150 295
<< nmos >>
rect -10 -300 5 -200
<< pmos >>
rect -10 -50 5 150
<< ndiff >>
rect -55 -210 -10 -200
rect -55 -295 -45 -210
rect -25 -295 -10 -210
rect -55 -300 -10 -295
rect 5 -210 50 -200
rect 5 -295 20 -210
rect 40 -295 50 -210
rect 5 -300 50 -295
<< pdiff >>
rect -55 140 -10 150
rect -55 -40 -45 140
rect -25 -40 -10 140
rect -55 -50 -10 -40
rect 5 140 50 150
rect 5 -40 20 140
rect 40 -40 50 140
rect 5 -50 50 -40
<< ndiffc >>
rect -45 -295 -25 -210
rect 20 -295 40 -210
<< pdiffc >>
rect -45 -40 -25 140
rect 20 -40 40 140
<< psubdiff >>
rect -60 -350 50 -340
rect -60 -385 -40 -350
rect 35 -385 50 -350
rect -60 -395 50 -385
<< nsubdiff >>
rect -60 220 55 230
rect -60 195 -40 220
rect 40 195 55 220
rect -60 185 55 195
<< psubdiffcont >>
rect -40 -385 35 -350
<< nsubdiffcont >>
rect -40 195 40 220
<< poly >>
rect -10 150 5 175
rect -10 -120 5 -50
rect -65 -130 5 -120
rect -65 -160 -50 -130
rect -25 -160 5 -130
rect -65 -170 5 -160
rect 30 -130 75 -120
rect 30 -160 40 -130
rect 65 -160 75 -130
rect 30 -170 75 -160
rect -10 -200 5 -170
rect -10 -315 5 -300
<< polycont >>
rect -50 -160 -25 -130
rect 40 -160 65 -130
<< locali >>
rect -55 220 50 225
rect -55 195 -40 220
rect 40 195 50 220
rect -55 190 50 195
rect -55 140 -15 190
rect -55 -40 -45 140
rect -25 -40 -15 140
rect -55 -45 -15 -40
rect 10 140 50 145
rect 10 -40 20 140
rect 40 -40 50 140
rect 10 -120 50 -40
rect -60 -130 -15 -120
rect -60 -160 -50 -130
rect -25 -160 -15 -130
rect -60 -170 -15 -160
rect 10 -130 75 -120
rect 10 -160 40 -130
rect 65 -160 75 -130
rect 10 -170 75 -160
rect -55 -210 -15 -205
rect -55 -295 -45 -210
rect -25 -295 -15 -210
rect 10 -210 50 -170
rect 10 -295 20 -210
rect 40 -295 50 -210
rect -55 -345 -15 -295
rect -55 -350 45 -345
rect -55 -385 -40 -350
rect 35 -385 45 -350
rect -55 -390 45 -385
<< viali >>
rect -25 195 25 220
rect -50 -160 -25 -130
rect 40 -160 65 -130
rect -25 -380 25 -355
<< metal1 >>
rect -160 220 165 235
rect -160 195 -25 220
rect 25 195 165 220
rect -160 180 165 195
rect -170 -130 -15 -120
rect -170 -160 -50 -130
rect -25 -160 -15 -130
rect -170 -170 -15 -160
rect 10 -130 140 -120
rect 10 -160 40 -130
rect 65 -160 140 -130
rect 10 -170 140 -160
rect -165 -355 160 -340
rect -165 -380 -25 -355
rect 25 -380 160 -355
rect -165 -395 160 -380
<< labels >>
rlabel metal1 105 195 125 215 1 VCC
rlabel metal1 90 -155 110 -135 1 Y
rlabel metal1 -155 -165 -135 -145 1 A
rlabel metal1 115 -380 135 -360 1 VSS
<< end >>
